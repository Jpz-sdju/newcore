module ifu (
    input backend_final_flush,
    babalala.....
);
    
endmodule