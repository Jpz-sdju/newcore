`define WORD_WIDTH 32
`define CACHELINE_SIZE 64 //byte
