`define WORD_WIDTH 32
`define xxx::??