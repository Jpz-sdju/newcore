module frontend (
    what?
);
    
endmodule