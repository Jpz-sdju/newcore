module dff #(
    parameter WIDTH=1
) (
    input [WIDTH-1:0] din,
    
);
    
endmodule